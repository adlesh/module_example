module int_stuff

import int_add
import int_swap
