module int_add

pub const (
        constant = 4
)
